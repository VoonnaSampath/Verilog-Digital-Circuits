module or4 (output y, input a, input b, input c, input d);
  or (y, a, b, c, d);
endmodule