module xor4 (output y, input a, input b, input c, input d);
  xor (y, a, b, c, d);
endmodule