module and4 (output y, input a, input b, input c, input d);
  and (y, a, b, c, d);
endmodule